interface dff_interface();
    logic din;
    logic clk;
    logic rst;
    logic dout;
  endinterface